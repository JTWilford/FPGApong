//////////////////////////////////////////////////////////////////////////////////
// Author:			Justin Wilford
// Create Date:		03/17/2019 
// File Name:		generate_pwm.v
// Description: 
//		Generates a PWM signal based on switch inputs.
//
// Revision: 		1.0
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module display_gandhi (
	input clk,
	input reset,
	//input sys_clk,
	input [10:0] ObjectX,		//Object's origin X Coordinate
	input [9:0] ObjectY,		//Object's origin Y Coordinate
	
	input [9:0] PollX,			//Position to Poll X Coordinate
	input [8:0] PollY,			//Position to Poll Y Coordinate
	
	output Hit,					//If HIGH, Then Poll Falls Within Object Bounds. Otherwise, LOW
	output Hit2
	);
	
	reg [9:0] TransformedPollX;
	reg [8:0] TransformedPollY;
	
	reg [99:0] GandhiMatrix [99:0];
	
	reg hit_out;
	reg hit2_out;
	
	//Get the ADC value from JPorts
	always @ (posedge clk)
	begin
		if(reset)
		begin
			hit_out <= 1'b0;
			hit2_out <= 1'b0;
			/*
			GandhiMatrix[0] <= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[1] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[2] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[3] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[4] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[5] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[6] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[7]  	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[8]  	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[9]  	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[10] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[11] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[12] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[13] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[14] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[15] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[16] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[17] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[18] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[19] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[20] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[21] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[22] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[23] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[24] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[25] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[26] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[27] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[28] 	<= 200'b00000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[29] 	<= 200'b00000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[30] 	<= 200'b00000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[31] 	<= 200'b00000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[32] 	<= 200'b00000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[33] 	<= 200'b00000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[34] 	<= 200'b00000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[35] 	<= 200'b00000000000000000000000000000000000000001100111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[36] 	<= 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[37] 	<= 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[38] 	<= 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[39] 	<= 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[40] 	<= 200'b00000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[41] 	<= 200'b00000000000000000000000000000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[42] 	<= 200'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[43] 	<= 200'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[44] 	<= 200'b00000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[45] 	<= 200'b00000000000000000000000000000000000000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[46] 	<= 200'b00000000000000000000000000000000000000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[47] 	<= 200'b00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[48] 	<= 200'b00000000000000000000000000000000000000000001111011111111111111111111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[49] 	<= 200'b00000000000000000000000000000000000000000001111001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[50] 	<= 200'b00000000000000000000000000000000000000000000111001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[51] 	<= 200'b00000000000000000000000000000000000000000000111001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[52] 	<= 200'b00000000000000000000000000000000000000000000111001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[53] 	<= 200'b00000000000000000000000000000000000000000000111001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[54] 	<= 200'b00000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[55] 	<= 200'b00000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[56] 	<= 200'b00000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[57] 	<= 200'b00000000000000000000000000000000000000000001111111111111111101111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[58] 	<= 200'b00000000000000000000000000000000000000000011111111000100000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[59] 	<= 200'b00000000000000000000000000000000000000000011111110000000000000000000000011111100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[60] 	<= 200'b00000000000000000000000000000000000000000011111100000000000000000000000011111000000011110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[61] 	<= 200'b00000000000000000000000000000000000000000011111000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[62] 	<= 200'b00000000000000000000000000000000000000000011111000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[63] 	<= 200'b00000000000000000000000000000000000000000011110000001111111000000000000001110000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[64] 	<= 200'b00000000000000000000000000000000000000000011100000001111111000000000000000100000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[65] 	<= 200'b00000000000000000000000000000000000000000011000000000000000000000000010000011100000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[66] 	<= 200'b00000000000000000000000000000000000000000011100000000000000001000000011000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[67] 	<= 200'b00000000000000000000000000000000000000000010000000000000000001100000110000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[68] 	<= 200'b00000000000000000000000000000000000000000000000000000010000001100000100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[69] 	<= 200'b00000000000000000000000000000000010000000000000000000011000000000000100001111110000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[70] 	<= 200'b00000000000000000000000000000000011111000011000000000011001000000000111001111111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[71] 	<= 200'b00000000000000000000000000000000011111100011100000000000000000000000011001111111000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[72] 	<= 200'b00000000000000000000000000000001111111110011000000000000000000000011110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[73] 	<= 200'b00000000000000000000000000000001111111110011100000000000000000000111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[74] 	<= 200'b00000000000000000000000000000001111111110011100000000000000000011111110011111111000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[75] 	<= 200'b00000000000000000000000000000001111111111011100000000000001111111111110111111111000000000000100001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[76] 	<= 200'b00000000000000000000000000000001111111111111110000111111111111111111100111111111000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[77] 	<= 200'b00000000000000000000000000000001111111111111100001111111111111111111111111111111000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[78] 	<= 200'b00000000000000000000000000000001111111111001111111111111111111111111111111111111000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[79] 	<= 200'b00000000000000000000000000000001111111111100111111111111111111111111111111111111100000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[80] 	<= 200'b00000000000000000000000000000001111111111110111111111111111111111111111111111111100000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[81] 	<= 200'b00000000000000000000000000000000111111111110111111111111111111111111111111111111110000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[82] 	<= 200'b00000000000000000000000000000000111111111111111111111111111111111111111111111111111000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[83] 	<= 200'b00000000000000000000000000000000011111111111011111111111111111111111111111111111111000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[84] 	<= 200'b00000000000000000000000000000000011111111111011111111111111111111111111111111111111000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[85] 	<= 200'b00000000000000000000000000000000011111111111011111111111111111111111111111111111111000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[86] 	<= 200'b00000000000000000000000000000000001111111111101111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[87] 	<= 200'b00000000000000000000000000000000001111111111101111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[88] 	<= 200'b00000000000000000000000000000000001111111111101111111111111111111111110011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[89] 	<= 200'b00000000000000000000000000000000000111111111110011111111111111110111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[90] 	<= 200'b00000000000000000000000000000000000111111111110011111111111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[91] 	<= 200'b00000000000000000000000000000000000111111111100011111111111110000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[92] 	<= 200'b00000000000000000000000000000000000111111111110000111111111110000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[93] 	<= 200'b00000000000000000000000000000000000011111111110000111111111100001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[94] 	<= 200'b00000000000000000000000000000000000011111111111000011111111000001101111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[95] 	<= 200'b00000000000000000000000000000000000011111111111100000111000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[96] 	<= 200'b00000000000000000000000000000000000001111111111100000101100000001111111111111111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[97] 	<= 200'b00000000000000000000000000000000000001111111111100000000000000101111100111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[98] 	<= 200'b00000000000000000000000000000000000000111111111100000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[99] 	<= 200'b00000000000000000000000000000000000000011111111000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[100]	<= 200'b00000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[101]	<= 200'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[102]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[103]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[104]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[105]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[106]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[107]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[108]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[109]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[110]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[111]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[112]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[113]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[114]	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000011111001001111001000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[115] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[116] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[117] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000011111111111001000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[118] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000001111111111001000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[119] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[120] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[121] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[122] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[123] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[124] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[125] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000110000011000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[126] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000011000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[127] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000111100000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[128] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111101011100000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[129] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111011100100000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[130] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111100100000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[131] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111101111100000111000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[132] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000101100000111111000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[133] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011000001110000011111000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[134] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011100001110000011111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[135] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011100000001000001111000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[136] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011110000001110000111000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[137] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011110000000110000011000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[138] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000011110000000001000011000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[139] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111000000001000001000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[140] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[141] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[142] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111110000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[143] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111000000000110001011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[144] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111110000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[145] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[146] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[147] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111111100011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[148] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[149] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[150] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[151] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111110111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[152] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111111111111100000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[153] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111111000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[154] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111110000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[155] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111110000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[156] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[157] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[158] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[159] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[160] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000111100000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[161] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000111110000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[162] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000011111100000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[163] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000111100000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[164] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[165] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[166] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[167] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[168] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[169] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[170] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111101000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[171] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111100000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[172] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[173] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111111000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[174] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000011000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[175] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000010000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[176] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000110000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[177] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111110000111000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[178] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111100000111000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[179] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111100001111000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[180] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111100001110000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[181] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111000001000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[182] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111000001000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[183] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111111000001100000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[184] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111110000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[185] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[186] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[187] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111110000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[188] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[189] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[190] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111100000000000110000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[191] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111100000000000110000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[192] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111100000000000100000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[193] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000001111000000011000100000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[194] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000000011000100000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[195] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000001001000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[196] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000111000001111000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[197] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000110000001111000000000001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[198] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000110000001111000000001001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[199] 	<= 200'b00000000000000000000000000000000000000000000000000000000000000000110000001110000000001111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			*/
			GandhiMatrix[0] 	<= 100'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[1] 	<= 100'b0000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000;
			GandhiMatrix[2] 	<= 100'b0000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000;
			GandhiMatrix[3] 	<= 100'b0000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000;
			GandhiMatrix[4] 	<= 100'b0000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[5] 	<= 100'b0000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[6] 	<= 100'b0000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[7] 	<= 100'b0000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[8] 	<= 100'b0000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[9] 	<= 100'b0000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[10] 	<= 100'b0000000000000110011111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[11] 	<= 100'b0000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000;
			GandhiMatrix[12] 	<= 100'b0000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[13] 	<= 100'b0000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[14] 	<= 100'b0000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[15] 	<= 100'b0000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[16] 	<= 100'b0000000000000011111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[17] 	<= 100'b0000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[18] 	<= 100'b0000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[19] 	<= 100'b0000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[20] 	<= 100'b0000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000;
			GandhiMatrix[21] 	<= 100'b0000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000;
			GandhiMatrix[22] 	<= 100'b0000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrix[23] 	<= 100'b0000000000000000111101111111111111111111111111111111111111111111010000000000000000000000000000000000;
			GandhiMatrix[24] 	<= 100'b0000000000000000111100111111111111111111111111111111111111111111111000000000000000000000000000000000;
			GandhiMatrix[25] 	<= 100'b0000000000000000011100111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrix[26] 	<= 100'b0000000000000000011100111111111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrix[27] 	<= 100'b0000000000000000011100111111111111111111111111111111111111110000000000000000000000000000000000000000;
			GandhiMatrix[28] 	<= 100'b0000000000000000011100111111111111111111111111111111111111100000000000000000000000000000000000000000;
			GandhiMatrix[29] 	<= 100'b0000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000;
			GandhiMatrix[30] 	<= 100'b0000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[31] 	<= 100'b0000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000;
			GandhiMatrix[32] 	<= 100'b0000000000000000111111111111111110111111111111111111110000000000000000000000000000000000000000000000;
			GandhiMatrix[33] 	<= 100'b0000000000000001111111100010000000000001111111111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[34] 	<= 100'b0000000000000001111111000000000000000000000001111110000000111111000000000000000000000000000000000000;
			GandhiMatrix[35] 	<= 100'b0000000000000001111110000000000000000000000001111100000001111011000000000000000000000000000000000000;
			GandhiMatrix[36] 	<= 100'b0000000000000001111100000000000000000000000000111110000000000000000000000000000000000000000000000000;
			GandhiMatrix[37] 	<= 100'b0000000000000001111100000000000000000000000000111100000000000000000000000000000000000000000000000000;
			GandhiMatrix[38] 	<= 100'b0000000000000001111000000111111100000000000000111000000000000000110000000000000000000000000000000000;
			GandhiMatrix[39] 	<= 100'b0000000000000001110000000111111100000000000000010000000000000001111000000000000000000000000000000000;
			GandhiMatrix[40] 	<= 100'b0000000000000001100000000000000000000000001000001110000000000001100000000000000000000000000000000000;
			GandhiMatrix[41] 	<= 100'b0000000000000001110000000000000000100000001100011111000000000000000000000000000000000000000000000000;
			GandhiMatrix[42] 	<= 100'b0000000000000001000000000000000000110000011000011111000000000000000000000000000000000000000000000000;
			GandhiMatrix[43] 	<= 100'b0000000000000000000000000001000000110000010000011111000000000000000000000000000000000000000000000000;
			GandhiMatrix[44] 	<= 100'b0000001000000000000000000001100000000000010000111111000000000001000000000000000000000000000000000000;
			GandhiMatrix[45] 	<= 100'b0000001111100001100000000001100100000000011100111111100000000001100000000000000000000000000000000000;
			GandhiMatrix[46] 	<= 100'b0000001111110001110000000000000000000000001100111111100000000000001111110000000000000000000000000000;
			GandhiMatrix[47] 	<= 100'b0000111111111001100000000000000000000001111000111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[48] 	<= 100'b0000111111111001110000000000000000000011111000111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[49] 	<= 100'b0000111111111001110000000000000000001111111001111111100000000000000000011111100000000000000000000000;
			GandhiMatrix[50] 	<= 100'b0000111111111101110000000000000111111111111011111111100000000000010000111111100000000000000000000000;
			GandhiMatrix[51] 	<= 100'b0000111111111111111000011111111111111111110011111111100000000000000111111111110000000000000000000000;
			GandhiMatrix[52] 	<= 100'b0000111111111111110000111111111111111111111111111111100000000000001111111111110000000000000000000000;
			GandhiMatrix[53] 	<= 100'b0000111111111100111111111111111111111111111111111111100000000000011111111111110000000000000000000000;
			GandhiMatrix[54] 	<= 100'b0000111111111110011111111111111111111111111111111111110000000000111111111111110000000000000000000000;
			GandhiMatrix[55] 	<= 100'b0000111111111111011111111111111111111111111111111111110000000000001111111111110000000000000000000000;
			GandhiMatrix[56] 	<= 100'b0000011111111111011111111111111111111111111111111111111000000000000111111111110000000000000000000000;
			GandhiMatrix[57] 	<= 100'b0000011111111111111111111111111111111111111111111111111100000000000011111111110000000000000000000000;
			GandhiMatrix[58] 	<= 100'b0000001111111111101111111111111111111111111111111111111100000000000001111111110000000000000000000000;
			GandhiMatrix[59] 	<= 100'b0000001111111111101111111111111111111111111111111111111100000000000000011111110000000000000000000000;
			GandhiMatrix[60] 	<= 100'b0000001111111111101111111111111111111111111111111111111100000000000000001111100000000000000000000000;
			GandhiMatrix[61] 	<= 100'b0000000111111111110111111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[62] 	<= 100'b0000000111111111110111111111111111111111111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[63] 	<= 100'b0000000111111111110111111111111111111111111001111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[64] 	<= 100'b0000000011111111111001111111111111111011100000001111111000000000000000000000000000000000000000000000;
			GandhiMatrix[65] 	<= 100'b0000000011111111111001111111111111100011111000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[66] 	<= 100'b0000000011111111110001111111111111000001111111111000000000000000000000000000000000000000000000000000;
			GandhiMatrix[67] 	<= 100'b0000000011111111111000011111111111000011111111111110000000000000000000000000000000000000000000000000;
			GandhiMatrix[68] 	<= 100'b0000000001111111111000011111111110000111111111111111100000000000000000000000000000000000000000000000;
			GandhiMatrix[69] 	<= 100'b0000000001111111111100001111111100000110111111111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[70] 	<= 100'b0000000001111111111110000011100000001111111111111111111000000000000000000000000000000000000000000000;
			GandhiMatrix[71] 	<= 100'b0000000000111111111110000010110000000111111111111111100011000000000000000000000000000000000000000000;
			GandhiMatrix[72] 	<= 100'b0000000000111111111110000000000000010111110011111111111110000000000000000000000000000000000000000000;
			GandhiMatrix[73] 	<= 100'b0000000000011111111110000000000000000000000001111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[74] 	<= 100'b0000000000001111111100000000000000000000000001111111111100000000000000000000000000000000000000000000;
			GandhiMatrix[75]	<= 100'b0000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[76]	<= 100'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[77]	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrix[78]	<= 100'b0000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000;
			GandhiMatrix[79]	<= 100'b0000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000;
			GandhiMatrix[80]	<= 100'b0000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000;
			GandhiMatrix[81]	<= 100'b0000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000;
			GandhiMatrix[82]	<= 100'b0000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000100000000;
			GandhiMatrix[83]	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
			GandhiMatrix[84]	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000;
			GandhiMatrix[85]	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000;
			GandhiMatrix[86]	<= 100'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011111000000;
			GandhiMatrix[87]	<= 100'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000000011111110000;
			GandhiMatrix[88]	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000;
			GandhiMatrix[89]	<= 100'b0000000000000000000000000000000000000000000001111100100111100100000000000000000000000000111111111000;
			GandhiMatrix[90] 	<= 100'b0000000000000000000000000000000000000000000000111111111111100000000000000000000000000001111111111000;
			GandhiMatrix[91] 	<= 100'b0000000000000000000000000000000000000000000000011111111111100000000000000000000000000001111111111000;
			GandhiMatrix[92] 	<= 100'b0000000000000000000000000000000000000000000000001111111111100100000000000000000000000011111111111000;
			GandhiMatrix[93] 	<= 100'b0000000000000000000000000000000000000000000000000111111111100100000000000000000000000011111111111000;
			GandhiMatrix[94] 	<= 100'b0000000000000000000000000000000000000000000000000011100111000000000000000000000000000111111111111000;
			GandhiMatrix[95] 	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000;
			GandhiMatrix[96] 	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000;
			GandhiMatrix[97] 	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000;
			GandhiMatrix[98] 	<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000;
			GandhiMatrix[99] 	<= 100'b0000000000000000000000000000000000000011000000000000000000000000000000000000000000111111111111100000;

		end
		else
		begin
			
			//Check if poll falls within the bounds of this object
			if((ObjectX <= PollX & PollX < ObjectX+100)&(ObjectY <= PollY & PollY < ObjectY+100))
				begin
					//Transform the polling coords
					TransformedPollX = PollX - ObjectX;
					TransformedPollY = PollY - ObjectY;
					
					hit_out <= GandhiMatrix[TransformedPollY][TransformedPollX];
					hit2_out <= ~GandhiMatrix[TransformedPollY][TransformedPollX];
				end
			else
				begin
				hit_out <= 1'b0;
				hit2_out <= 1'b0;
				end
		end
	end
	
	assign Hit = hit_out;
	assign Hit2 = hit2_out;

endmodule