//////////////////////////////////////////////////////////////////////////////////
// Author:			Justin Wilford
// Create Date:		04/17/2019 
// File Name:		display_gandhi.v
// Description: 
//		Displays a 100px by 100px monochromatic image of Professor Gandhi Puvvada.
//
// Revision: 		1.1
// Additional Comments:  Was originally 200px by 200px, but ISE ran out of memory while synthesizing.
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module display_gandhi (
	input clk,
	input reset,
	//input sys_clk,
	input [10:0] ObjectX,		//Object's origin X Coordinate
	input [9:0] ObjectY,		//Object's origin Y Coordinate
	
	input [9:0] PollX,			//Position to Poll X Coordinate
	input [8:0] PollY,			//Position to Poll Y Coordinate
	
	output Hit,					//If HIGH, Then Poll Falls Within Object Bounds. Otherwise, LOW
	output Hit2
	);
	
	reg [9:0] TransformedPollX;
	reg [8:0] TransformedPollY;
	
	reg [99:0] GandhiMatrixReverse [99:0];
	reg [99:0] GandhiMatrixNormal [99:0];
	
	reg hit_out;
	reg hit2_out;
	
	//Get the ADC value from JPorts
	always @ (posedge clk)
	begin
		if(reset)
		begin
			hit_out <= 1'b0;
			hit2_out <= 1'b0;
			
			GandhiMatrixReverse[0] 		<= 100'b0000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000;
			GandhiMatrixReverse[1] 		<= 100'b0000000000000000000000000000000000000000001111000000000111111111110000000000000000000000000000000000;
			GandhiMatrixReverse[2] 		<= 100'b0000000000000000000000000000000000000001111111000000000001111111111100000000000000000000000000000000;
			GandhiMatrixReverse[3] 		<= 100'b0000000000000000000000000000000000001111110000000000000000011111111110000000000000000000000000000000;
			GandhiMatrixReverse[4] 		<= 100'b0000000000000000000000000000000001111100000000000000000000000011111111000000000000000000000000000000;
			GandhiMatrixReverse[5] 		<= 100'b0000000000000000000000000000001111111000000000000000000000000001111111100000000000000000000000000000;
			GandhiMatrixReverse[6] 		<= 100'b0000000000000000000001100000111100000000000000000000000000000000111111100000000000000000000000000000;
			GandhiMatrixReverse[7] 		<= 100'b0000000000000000000011000111111000000000001110000000000000000000111111100000000000000000000000000000;
			GandhiMatrixReverse[8] 		<= 100'b0000000000000000000011100111100000000000011111111000000000000000111111100000000000000000000000000000;
			GandhiMatrixReverse[9] 		<= 100'b0000000000000000000111011111000000001100011111110000000000000001111111110000000000000000000000000000;
			GandhiMatrixReverse[10] 	<= 100'b0000000000000000001111111100000000111111110111111000000000000000111111110000000000000000000000000000;
			GandhiMatrixReverse[11] 	<= 100'b0000000000000000001011100000000001111111111000011000000000000000111111110000000000000000000000000000;
			GandhiMatrixReverse[12] 	<= 100'b0000000000000000010001000000000111111111111111110000000000000001111111110000000000000000000000000000;
			GandhiMatrixReverse[13] 	<= 100'b0000000000000000011100000000001111111111111111110000000000000001111111111000000000000000000000000000;
			GandhiMatrixReverse[14] 	<= 100'b0000001000000000001100000000001111111111111111110000000000000000001111111000000000000000000000000000;
			GandhiMatrixReverse[15] 	<= 100'b0000001000000000001111100000011111111111111111111000000000000000011111111100000000000000000000000000;
			GandhiMatrixReverse[16] 	<= 100'b0000000000000000011111100000011111111111111110111100000000000000011111111100000000000000000000000000;
			GandhiMatrixReverse[17] 	<= 100'b0000000000000000001111100000001111111111111110011100000000000000011111111100000000000000000000000000;
			GandhiMatrixReverse[18] 	<= 100'b0000000000010000001111100000011111111111111111111100000000000000011111111100000000000000000000000000;
			GandhiMatrixReverse[19] 	<= 100'b0000000000010100001111000000001111111111111111111000000000000000011111111100000000000000000000000000;
			GandhiMatrixReverse[20] 	<= 100'b0000000000000100001111000000001111111111111111110110000000000000001111111110000000000000000000000000;
			GandhiMatrixReverse[21] 	<= 100'b0000000000001110001111000000001111111111111111110111100000000000000111111110000000000000000000000000;
			GandhiMatrixReverse[22] 	<= 100'b0000000000111110101100000000001111111111111110111111100000000000000011111110000000000000000000000000;
			GandhiMatrixReverse[23] 	<= 100'b0000000000011100100100000000000111111111011100000011100000000000000001111110000000000000000000000000;
			GandhiMatrixReverse[24] 	<= 100'b0000000000011101100110000000000000000000000000000001100000000000000000011111000000000000000000000000;
			GandhiMatrixReverse[25] 	<= 100'b0000000000001100100110000000000000000000000000000001100000000000000000000111000000000000000000000000;
			GandhiMatrixReverse[26] 	<= 100'b0000000000011100100110000000000000111110000000000001100000000000000000000111000000000000000000000000;
			GandhiMatrixReverse[27] 	<= 100'b0000000000011100100110000000000001111111110000000011111100000000000000011111000000000000000000000000;
			GandhiMatrixReverse[28] 	<= 100'b0000000000111100101110000000000000011111110000000011111111101100000001111100000000000000000000000000;
			GandhiMatrixReverse[29] 	<= 100'b0000000000111110001110000000000000011111111111000011111111110000001111100000000000000000000000000000;
			GandhiMatrixReverse[30] 	<= 100'b0000000000010110011110000000001111111111111111100011111111110000110000000000000000000000000000000000;
			GandhiMatrixReverse[31] 	<= 100'b0100000000000010011110000000011111111111111111110011111111100001100000000000000000000000000000000000;
			GandhiMatrixReverse[32] 	<= 100'b0100000000000010001110000000011111111111111111110011111111000110000000000000000000000000000000000000;
			GandhiMatrixReverse[33] 	<= 100'b0000000000000010000011100000011111111111111111111011111110001100000001111000000000000000000000000000;
			GandhiMatrixReverse[34] 	<= 100'b0000000000000010000101100000001110000000000011100011100000011000000011100000000000000000000000000000;
			GandhiMatrixReverse[35] 	<= 100'b0000000000000101000100000000000001110011111000000001100000110000011111111100000000000000000000000000;
			GandhiMatrixReverse[36] 	<= 100'b0000000000000111000100111001111110000000111110000001100011100010011001011000000000000000000000000000;
			GandhiMatrixReverse[37] 	<= 100'b0000000000001111000101111001000000000000000011111001100011101111001001110000000000000000000000000000;
			GandhiMatrixReverse[38] 	<= 100'b0000000000001110000011110010000000000000000000001101110011001000111111000000110000000000000000000000;
			GandhiMatrixReverse[39] 	<= 100'b0000000000000000000010000111111110101111100000000001110011001111111110100000110000000000000000000000;
			GandhiMatrixReverse[40] 	<= 100'b0000000000000000000010001100110111111110001111100000110110001111001111110000111000000000000000000000;
			GandhiMatrixReverse[41] 	<= 100'b0000000000000000000010011001111111000111000011100011001000000001111101100111110000000000000000000000;
			GandhiMatrixReverse[42] 	<= 100'b0000000000000000000100101111111111110001000011100001000001000001111000001111100000000000000000000000;
			GandhiMatrixReverse[43] 	<= 100'b0000000000000000000010011111111110000000110011000001111001000000111001111111000000000000000000000000;
			GandhiMatrixReverse[44] 	<= 100'b0000000000000000000101111111000110000000011111001001100001100000011111111100000000000000000000000000;
			GandhiMatrixReverse[45] 	<= 100'b0000000001111000000100001111000101000010011111011000011100100000011111111111000001111100000000000000;
			GandhiMatrixReverse[46] 	<= 100'b0000000011001111011100000110000110101111111011011010111000100000011000111111111111111100000000000000;
			GandhiMatrixReverse[47] 	<= 100'b0000000011000000011100100100000100010111100010000111111000100000001100000011001111011000000000000000;
			GandhiMatrixReverse[48] 	<= 100'b0000000011100000011100000000000111011111001100000111111100100000111100000000001111111110000000000000;
			GandhiMatrixReverse[49] 	<= 100'b0000000010000000001010010001101111111111111000000011111100110000001110000111111111111111000000000000;
			GandhiMatrixReverse[50] 	<= 100'b0000000011101111001111010011111111001111110000001001111100110000000000000111110000011111000000000000;
			GandhiMatrixReverse[51] 	<= 100'b0000000011101111100111010011111111111110000011100101111100110010000111111110000000001111000000000000;
			GandhiMatrixReverse[52] 	<= 100'b0000000001101111110100001011100111000000000000000000111100110001111110000000000000000111000000000000;
			GandhiMatrixReverse[53] 	<= 100'b0000000001111111110000001111000000011110000000000000011100111001111111000000000000000111000000000000;
			GandhiMatrixReverse[54] 	<= 100'b0000000001111111110000000010000000011111111100001100011100111000111111000000001100001111100000000000;
			GandhiMatrixReverse[55] 	<= 100'b0000000001111111110010000001100000000000000000000000011110010000111110000000000000001111000000000000;
			GandhiMatrixReverse[56] 	<= 100'b0000000011111111100010000000000000000000000000111110011110010000011110000000000000001111000000000000;
			GandhiMatrixReverse[57] 	<= 100'b0000000001111111100000000000110011000000000001110000011111011000111011000000000000001111000000000000;
			GandhiMatrixReverse[58] 	<= 100'b0000000000111111000000000001111111111111110000000000011111001101111100100000000000001111000000000000;
			GandhiMatrixReverse[59] 	<= 100'b0000000001111111001100000001111111111111110111000000001111000101101100011000000000001111000000000000;
			GandhiMatrixReverse[60] 	<= 100'b0000000000011110001110000011111111111111111110000000001110000110111110001100000000001110000000000000;
			GandhiMatrixReverse[61] 	<= 100'b0000000000111110001110000011111111111111111100000000011111000011111100000110000000001110000000000000;
			GandhiMatrixReverse[62] 	<= 100'b0000000000011111011110000111111111111111111000011000011111100011100000000011000000001110000000000000;
			GandhiMatrixReverse[63] 	<= 100'b0000000000011111011110000001111111111111110000111000011111100011000000000001110000111100000000000000;
			GandhiMatrixReverse[64] 	<= 100'b0000000000001111001110000000111111111111000000000000111111110010000000000000111111111100000000000000;
			GandhiMatrixReverse[65] 	<= 100'b0000000000001111100110000000111111111110000000000000011111100110000000000000001111111100000000000000;
			GandhiMatrixReverse[66] 	<= 100'b0000000000001111100000000000111111111110000000001111000000001100000000000000011001111000000000000000;
			GandhiMatrixReverse[67] 	<= 100'b0000000000000111100000000000111111111100011000000111111000011000000011110000010001110000000000000000;
			GandhiMatrixReverse[68] 	<= 100'b0000000000000111111000000000000111111000111000000000000011100000000111111000010100111000000000000000;
			GandhiMatrixReverse[69] 	<= 100'b0000000000000111111110000100000011100001110000000000000001110011111111111000000000111000000000000000;
			GandhiMatrixReverse[70] 	<= 100'b0000000000000011111111000110000000000011110000000000000000111111111111111000000010111000000000000000;
			GandhiMatrixReverse[71] 	<= 100'b0000000000000011111111100011000000000011100000000000000000000001111111110000000011111000000000000000;
			GandhiMatrixReverse[72] 	<= 100'b0000000000000011111111110011000000000111100000000000000000000000111111110000000011111000000000000000;
			GandhiMatrixReverse[73] 	<= 100'b0000000000000011111111111101110000001101000000000000000000000000101111000000000011110000000000000000;
			GandhiMatrixReverse[74] 	<= 100'b0000000000000001111111111001111000001111000000000000000000000000111111000000000011110000000000000000;
			GandhiMatrixReverse[75]		<= 100'b0000000000000000111111111011111111011111011100000000000000000011111100000000000111110000000000000000;
			GandhiMatrixReverse[76]		<= 100'b0000000000000000111111110000111111111111111111100000000000000111101000000000000111100000000000000000;
			GandhiMatrixReverse[77]		<= 100'b0000000000000000010111101100111111111111100011111100000001111111100000000000000111100000000000000000;
			GandhiMatrixReverse[78]		<= 100'b0000000000000000001100011000111111111111000111111111111111111000000000000000000111000000000000000000;
			GandhiMatrixReverse[79]		<= 100'b0000000000000000000000000000011111111111101111111110111111000001111110000000000110000000000000001000;
			GandhiMatrixReverse[80]		<= 100'b0000000000000000000000000000011111111110111111111111111111111110000100000000000000000000000000001000;
			GandhiMatrixReverse[81]		<= 100'b0000000000000000000000000000011111111111111111111111100000000000000100000000000000000000000000001100;
			GandhiMatrixReverse[82]		<= 100'b0000000000000000000000000000001111111111111111111111100001100000011100000000000000000000000000001100;
			GandhiMatrixReverse[83]		<= 100'b0000000000000000000000000000000111111111111111111111100000000000011000000000000000000000000000011110;
			GandhiMatrixReverse[84]		<= 100'b0000000000000000000000000000000111111111111111011111110000000001110000000000000000000000000000010110;
			GandhiMatrixReverse[85]		<= 100'b0000000000000000000000000000000011111111111110000111111111011110000000000000000000000000000000000110;
			GandhiMatrixReverse[86]		<= 100'b0000000000000000000000000000000001111111111110000011111111110000000001111100000000000000000000100011;
			GandhiMatrixReverse[87]		<= 100'b0000000000000000000000000000000001111111111110000001111111111111100111111110000000000000000000100011;
			GandhiMatrixReverse[88]		<= 100'b0000000000000000000000000000000000111111111111100000111111111111111111111110000000000000000000000000;
			GandhiMatrixReverse[89]		<= 100'b0000000000000000000000000000000000011111111111110000110111111111111111111100000000000000000001000000;
			GandhiMatrixReverse[90] 	<= 100'b0000000000000000000000000000000000001111111111111000000001111111110111111100000000000000000000000000;
			GandhiMatrixReverse[91] 	<= 100'b0000000000000000000000000000000000000111111111111100000000000000000011111100000000000000000010000000;
			GandhiMatrixReverse[92] 	<= 100'b0000000000000000000000000000000000000001111111111100000000000000000011111000000000000000000011101110;
			GandhiMatrixReverse[93] 	<= 100'b0000000000000000000000000000000000000000111111111110000000000000000011110000000000000000000011111110;
			GandhiMatrixReverse[94] 	<= 100'b0000000000000000000000000000000000000000011111111111000000000000000011110000000000000000000111111110;
			GandhiMatrixReverse[95] 	<= 100'b0000000000000000000000000000000000000000011111111111100000000000000111100000000000000000000111111111;
			GandhiMatrixReverse[96] 	<= 100'b0000000000000000000000000000000000000000011100111111111000000000001111000000000000000000001111111111;
			GandhiMatrixReverse[97] 	<= 100'b0000000000000000000000000000000000000000011111001111111000100001111110000000000000000000001111111111;
			GandhiMatrixReverse[98] 	<= 100'b0000000000000000000000000000000000000000011011101011111111111111111000000000000000000000011111111111;
			GandhiMatrixReverse[99] 	<= 100'b0000000000000000000000000000000000000000111011111110011111111110000000000000000000000000011111111111;
			
			GandhiMatrixNormal[0] 		<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrixNormal[1] 		<= 100'b0000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000;
			GandhiMatrixNormal[2] 		<= 100'b0000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000;
			GandhiMatrixNormal[3] 		<= 100'b0000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000;
			GandhiMatrixNormal[4] 		<= 100'b0000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000;
			GandhiMatrixNormal[5] 		<= 100'b0000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[6] 		<= 100'b0000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[7] 		<= 100'b0000000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[8] 		<= 100'b0000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[9] 		<= 100'b0000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[10] 		<= 100'b0000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[11] 		<= 100'b0000000000000000000100011111111111111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[12] 		<= 100'b0000000000000000001110111111111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[13] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[14] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000;
			GandhiMatrixNormal[15] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[16] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[17] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[18] 		<= 100'b0000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[19] 		<= 100'b0000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[20] 		<= 100'b0000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000000000000;
			GandhiMatrixNormal[21] 		<= 100'b0000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000;
			GandhiMatrixNormal[22] 		<= 100'b0000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000;
			GandhiMatrixNormal[23] 		<= 100'b0000000000000000000011111111111111111111111111111111111111111111111110000000000000000000000000000000;
			GandhiMatrixNormal[24] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000;
			GandhiMatrixNormal[25] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000;
			GandhiMatrixNormal[26] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000;
			GandhiMatrixNormal[27] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000;
			GandhiMatrixNormal[28] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000;
			GandhiMatrixNormal[29] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000;
			GandhiMatrixNormal[30] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[31] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[32] 		<= 100'b0000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000;
			GandhiMatrixNormal[33] 		<= 100'b0000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000;
			GandhiMatrixNormal[34] 		<= 100'b0000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000;
			GandhiMatrixNormal[35] 		<= 100'b0000000000000000000011111111111110000000000111111111111111000000000000000000000000000000000000000000;
			GandhiMatrixNormal[36] 		<= 100'b0000000000000000000011111110000000000000000001111111111100000001111110100000000000000000000000000000;
			GandhiMatrixNormal[37] 		<= 100'b0000000000000000000011111110000000000000000000000111111100000011110110000000000000000000000000000000;
			GandhiMatrixNormal[38] 		<= 100'b0000000000000000000011111100000000000000000000000011111100000111000000000000000000000000000000000000;
			GandhiMatrixNormal[39] 		<= 100'b0000000000000000000011111000000001010000000000000011111100000000000001000000000000000000000000000000;
			GandhiMatrixNormal[40] 		<= 100'b0000000000000000000011110000001111111000000000000011111000000000110011100000000000000000000000000000;
			GandhiMatrixNormal[41] 		<= 100'b0000000000000000000011100000001111111000000000011000110000000000000011111000000000000000000000000000;
			GandhiMatrixNormal[42] 		<= 100'b0000000000000000000011000000000000000000000000011000111110000000000111110000000000000000000000000000;
			GandhiMatrixNormal[43] 		<= 100'b0000000000000000000011100000000000000001000000111000111110000000000110000000000000000000000000000000;
			GandhiMatrixNormal[44] 		<= 100'b0000000000000000000010000000000000000001100000110001111110000000000000000000000000000000000000000000;
			GandhiMatrixNormal[45] 		<= 100'b0000000000000000000000000000000010000001100000100001111111000000000000000000000000000000000000000000;
			GandhiMatrixNormal[46] 		<= 100'b0000000000110000000000000000000111000000000000100001111111000000000111000000000000000000000000000000;
			GandhiMatrixNormal[47] 		<= 100'b0000000000111111100011000000000011101000000001111001111111000000000011111100110000000000000000000000;
			GandhiMatrixNormal[48] 		<= 100'b0000000000011111100011100000000000100000000011111001111111000000000011111111110000000000000000000000;
			GandhiMatrixNormal[49] 		<= 100'b0000000001111111110011100000000000000000000111111001111111000000000001111000000000000000000000000000;
			GandhiMatrixNormal[50] 		<= 100'b0000000001111111110011100000000000110000001111110011111111000000000000000000001111100000000000000000;
			GandhiMatrixNormal[51] 		<= 100'b0000000001111111111011100000000000000001111111111011111111000000000000000001111111110000000000000000;
			GandhiMatrixNormal[52] 		<= 100'b0000000001111111111011110000011000111111111111111111111111000000000001111111111111111000000000000000;
			GandhiMatrixNormal[53] 		<= 100'b0000000001111111111111110000111111111111111111111111111111000000000000111111111111111000000000000000;
			GandhiMatrixNormal[54] 		<= 100'b0000000001111111111111111101111111111111111111111111111111000000000000111111111111110000000000000000;
			GandhiMatrixNormal[55] 		<= 100'b0000000001111111111101111111111111111111111111111111111111100000000001111111111111110000000000000000;
			GandhiMatrixNormal[56] 		<= 100'b0000000001111111111101111111111111111111111111111111111111100000000001111111111111110000000000000000;
			GandhiMatrixNormal[57] 		<= 100'b0000000001111111111111111111111111111111111111111111111111100000000000111111111111110000000000000000;
			GandhiMatrixNormal[58] 		<= 100'b0000000000111111111111111111111111111111111111111111111111110000000000011111111111110000000000000000;
			GandhiMatrixNormal[59] 		<= 100'b0000000000111111111111111111111111111111111111111111111111111000010000000111111111110000000000000000;
			GandhiMatrixNormal[60] 		<= 100'b0000000000011111111111111111111111111111111111111111111111111000000000000011111111110000000000000000;
			GandhiMatrixNormal[61] 		<= 100'b0000000000011111111111111111111111111111111111111111111111111100000000000001111111110000000000000000;
			GandhiMatrixNormal[62] 		<= 100'b0000000000011111111111111111111111111111111111111111111111111100000000000000111111110000000000000000;
			GandhiMatrixNormal[63] 		<= 100'b0000000000001111111111111111111111111111111111111111111111111100000000000000001111000000000000000000;
			GandhiMatrixNormal[64] 		<= 100'b0000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000;
			GandhiMatrixNormal[65] 		<= 100'b0000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000;
			GandhiMatrixNormal[66] 		<= 100'b0000000000001111111111111111111111111111111111110000111111110000000000000000000000000000000000000000;
			GandhiMatrixNormal[67] 		<= 100'b0000000000000111111111111111111111111111100111111000000111100000000000000000000000000000000000000000;
			GandhiMatrixNormal[68] 		<= 100'b0000000000000111111111111111111111111111000111111111111100000000000000000000000000000000000000000000;
			GandhiMatrixNormal[69] 		<= 100'b0000000000000111111111111011111111111110001111111111111110000000000000000000000000000000000000000000;
			GandhiMatrixNormal[70] 		<= 100'b0000000000000011111111111001111111111100001111111111111111000000000000000000000000000000000000000000;
			GandhiMatrixNormal[71] 		<= 100'b0000000000000011111111111100111111111100011111111111111111111110000000000000000000000000000000000000;
			GandhiMatrixNormal[72] 		<= 100'b0000000000000011111111111100111111111000011111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[73] 		<= 100'b0000000000000011111111111110001111110000111111111111111111111111010000000000000000000000000000000000;
			GandhiMatrixNormal[74] 		<= 100'b0000000000000001111111111110000111110000111111111111111111111111000000000000000000000000000000000000;
			GandhiMatrixNormal[75]		<= 100'b0000000000000001111111111100000000100000100011111111111111111100000000000000000000000000000000000000;
			GandhiMatrixNormal[76]		<= 100'b0000000000000000011111111100000000000000000000011111111111111000000000000000000000000000000000000000;
			GandhiMatrixNormal[77]		<= 100'b0000000000000000001111110000000000000000000000000011111110000000000000000000000000000000000000000000;
			GandhiMatrixNormal[78]		<= 100'b0000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrixNormal[79]		<= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			GandhiMatrixNormal[80]		<= 100'b0000000000000000000000000000000000000001000000000000000000000001111000000000000000000000000000000000;
			GandhiMatrixNormal[81]		<= 100'b0000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000;
			GandhiMatrixNormal[82]		<= 100'b0000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[83]		<= 100'b0000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000;
			GandhiMatrixNormal[84]		<= 100'b0000000000000000000000000000000000000000000000100000001111111110000000000000000000000000000000001000;
			GandhiMatrixNormal[85]		<= 100'b0000000000000000000000000000000000000000000001111000000000100000000000000000000000000000000000011000;
			GandhiMatrixNormal[86]		<= 100'b0000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000011100;
			GandhiMatrixNormal[87]		<= 100'b0000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000011100;
			GandhiMatrixNormal[88]		<= 100'b0000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000111111;
			GandhiMatrixNormal[89]		<= 100'b0000000000000000000000000000000000000000000000001111001000000000000000000000000000000000000000111111;
			GandhiMatrixNormal[90] 		<= 100'b0000000000000000000000000000000000000000000000000111111110000000001000000000000000000000000001111111;
			GandhiMatrixNormal[91] 		<= 100'b0000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000001111111;
			GandhiMatrixNormal[92] 		<= 100'b0000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000011111111;
			GandhiMatrixNormal[93] 		<= 100'b0000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000011111111;
			GandhiMatrixNormal[94] 		<= 100'b0000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000111111111;
			GandhiMatrixNormal[95] 		<= 100'b0000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000111111111;
			GandhiMatrixNormal[96] 		<= 100'b0000000000000000000000000000000000000000000000000000000111111111110000000000000000000000001111111111;
			GandhiMatrixNormal[97] 		<= 100'b0000000000000000000000000000000000000000000000000000000111011110000000000000000000000000001111111111;
			GandhiMatrixNormal[98] 		<= 100'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000011111111111;
			GandhiMatrixNormal[99] 		<= 100'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000000011111111111;



		end
		else
		begin
			
			//Check if poll falls within the bounds of this object
			if((ObjectX <= PollX & PollX < ObjectX+100)&(ObjectY <= PollY & PollY < ObjectY+100))
				begin
					//Transform the polling coords
					TransformedPollX = PollX - ObjectX;
					TransformedPollY = PollY - ObjectY;
					
					case({GandhiMatrixNormal[TransformedPollY][TransformedPollX],GandhiMatrixReverse[TransformedPollY][TransformedPollX]})
						2'b00:
							begin
								hit_out <= 1'b0;
								hit2_out <= 1'b0;
							end
						2'b01:
							begin
								hit_out <= 1'b1;
								hit2_out <= 1'b0;
							end
						2'b10:
							begin
								hit_out <= 1'b0;
								hit2_out <= 1'b1;
							end
						2'b11:
							begin
								hit_out <= 1'b1;
								hit2_out <= 1'b1;
							end
					endcase
				end
			else
				begin
				hit_out <= 1'b0;
				hit2_out <= 1'b0;
				end
		end
	end
	
	assign Hit = hit_out;
	assign Hit2 = hit2_out;

endmodule